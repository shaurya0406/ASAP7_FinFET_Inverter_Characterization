** sch_path: /home/parallels/ASAP7_FinFET_Inverter_Characterization/Xschem_ASAP7/inverter_test.sch
**.subckt inverter_test
x1 vdd vin vout GND inverter
vdd vdd GND 0.7
vin vin GND PULSE(0 0.7 0p 10p 10p 20p 60p 2)
**** begin user architecture code



.control
run
set filetype=ascii
set appendwrite

echo "WPfet,WNfet,Vm,Id,Gain,NMH,NML,Gm,tpd,tRise,tFall,Fsw,Power,Rout" > results.csv
let wpfet = 6
foreach wpfet 14 13 12 11 10 9 8 7 6 5 4 3 2
	foreach wnfet 14 13 12 11 10 9 8 7 6 5 4 3 2
		alter n.x1.xpfet1.npmos_finfet nfin = $wpfet
      		alter n.x1.xnfet1.nnmos_finfet nfin = $wnfet
		show n.x1.xpfet1.npmos_finfet : nfin
      		show n.x1.xnfet1.nnmos_finfet : nfin

		dc vin 0 0.7 1m

		set brushwidth 3

		setplot dc
		*plot vin vout
		meas dc vm when vin=vout

		if $&dc.vm > 0.34
			if $&dc.vm < 0.36

				let id = abs(vdd#branch)
				meas dc id_max MAX id
				print id_max

				let gm = real(deriv(id, vin))
				meas dc gm_max MAX gm
				print gm_max

				let rout = abs(real(deriv(vout, id)))
				meas dc rout_max MAX rout
				print rout_max

				let gain = abs(deriv(vout))
				meas dc gain_max MAX gain
				let gain_scaled = (gain >= 1)*0.7
				*plot gain_scaled vout
				meas dc vil find vin when gain_scaled=0.7 cross=1
				meas dc vih find vin when gain_scaled=0.7 cross=last
				let vol = 0
				let voh = 0.7
				let nmh = voh-vih
				let nml = vil-vol
				print nmh
				print nml

				tran 0.02p 125p
				setplot tran

				*plot vin vout
				meas tran tin_rise50 when vin=0.35 RISE=2
				meas tran tout_fall50 when vout=0.35 FALL=2
				meas tran tin_fall50 when vin=0.35 FALL=2
				meas tran tout_rise50 when vout=0.35 RISE=2
				meas tran tout_rise10 when vout=0.07 RISE=2
				meas tran tout_rise90 when vout=0.63 RISE=2
				meas tran tout_fall10 when vout=0.07 FALL=2
				meas tran tout_fall90 when vout=0.63 FALL=2

				let tpHL = tout_fall50-tin_rise50
				let tpLH = tout_rise50-tin_fall50
				let tpd = (tpHL+tpLH)/2
				let tr = tout_rise90 - tout_rise10
				let tf = tout_fall10 - tout_fall90
				let fsw = 1/(tr+tf)
				let id_tran = vdd#branch
				*plot id*1000 vout
				meas tran id_integ integ id_tran from=60e-12 to=120e-12
				let power_int = id_integ*0.7
				let power = abs(power_int/60)

				print tpHL
				print tpLH
				print tpd
				print tr
				print tf
				print fsw
				print power


				echo "$wpfet,$wnfet,$&dc.vm,$&dc.id_max,$&dc.gain_max,$&dc.nmh,$&dc.nml,$&dc.gm_max,$&tran.tpd,$&tran.tr,$&tran.tf,$&tran.fsw,$&tran.power,$&dc.rout_max" >> results.csv
			end
		end
   	end
	*$&wpfet = $&wpfet-1
end


.endc
.save all
.end


**** end user architecture code
**.ends

* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/parallels/ASAP7_FinFET_Inverter_Characterization/Xschem_ASAP7/inverter.sym
** sch_path: /home/parallels/ASAP7_FinFET_Inverter_Characterization/Xschem_ASAP7/inverter.sch
.subckt inverter vdd vin vout gnd
*.ipin vin
*.ipin vdd
*.ipin gnd
*.opin vout
Xnfet1 vout vin gnd gnd asap_7nm_nfet l=7e-009 nfin=13
Xpfet1 vout vin vdd vout asap_7nm_pfet l=7e-009 nfin=14
.ends

.GLOBAL GND
**** begin user architecture code

.subckt asap_7nm_pfet S G D B l=7e-009 nfin=14
	npmos_finfet S G D B BSIMCMG_osdi_P l=7e-009 nfin=14
.ends asap_7nm_pfet

.model BSIMCMG_osdi_P BSIMCMG_va (
+ TYPE = 0

************************************************************
*                         general                          *
************************************************************
+version = 107             bulkmod = 1               igcmod  = 1               igbmod  = 0
+gidlmod = 1               iimod   = 0               geomod  = 1               rdsmod  = 0
+rgatemod= 0               rgeomod = 0               shmod   = 0               nqsmod  = 0
+coremod = 0               cgeomod = 0               capmod  = 0               tnom    = 25
+eot     = 1e-009          eotbox  = 1.4e-007        eotacc  = 3e-010          tfin    = 6.5e-009
+toxp    = 2.1e-009        nbody   = 1e+022          phig    = 4.9278          epsrox  = 3.9
+epsrsub = 11.9            easub   = 4.05            ni0sub  = 1.1e+016        bg0sub  = 1.17
+nc0sub  = 2.86e+025       nsd     = 2e+026          ngate   = 0               nseg    = 5
+l       = 2.1e-008        xl      = 1e-009          lint    = -2.5e-009       dlc     = 0
+dlbin   = 0               hfin    = 3.2e-008        deltaw  = 0               deltawcv= 0
+sdterm  = 0               epsrsp  = 3.9             nfin    = 1
+toxg    = 1.8e-009
************************************************************
*                            dc                            *
************************************************************
+cit     = 0               cdsc    = 0.003469        cdscd   = 0.001486        dvt0    = 0.05
+dvt1    = 0.36            phin    = 0.05            eta0    = 0.094           dsub    = 0.24
+k1rsce  = 0               lpe0    = 0               dvtshift= 0               qmfactor= 0
+etaqm   = 0.54            qm0     = 2.183e-012      pqm     = 0.66            u0      = 0.0237
+etamob  = 4               up      = 0               ua      = 1.133           eu      = 0.05
+ud      = 0.0105          ucs     = 0.2672          rdswmin = 0               rdsw    = 200
+wr      = 1               rswmin  = 0               rdwmin  = 0               rshs    = 0
+rshd    = 0               vsat    = 60000           deltavsat= 0.17            ksativ  = 1.592
+mexp    = 2.491           ptwg    = 25              pclm    = 0.01            pclmg   = 1
+pdibl1  = 800             pdibl2  = 0.005704        drout   = 4.97            pvag    = 200
+fpitch  = 2.7e-008        rth0    = 0.15            cth0    = 1.243e-006      wth0    = 2.6e-007
+lcdscd  = 0               lcdscdr = 0               lrdsw   = 1.3             lvsat   = 1441
************************************************************
*                         leakage                          *
************************************************************
+aigc    = 0.007           bigc    = 0.0015          cigc    = 1               dlcigs  = 5e-009
+dlcigd  = 5e-009          aigs    = 0.006           aigd    = 0.006           bigs    = 0.001944
+bigd    = 0.001944        cigs    = 1               cigd    = 1               poxedge = 1.152
+agidl   = 2e-012          agisl   = 2e-012          bgidl   = 1.5e+008        bgisl   = 1.5e+008
+egidl   = 1.142           egisl   = 1.142
************************************************************
*                            rf                            *
************************************************************
************************************************************
*                         junction                         *
************************************************************
************************************************************
*                       capacitance                        *
************************************************************
+cfs     = 0               cfd     = 0               cgso    = 1.6e-010        cgdo    = 1.6e-010
+cgsl    = 0               cgdl    = 0               ckappas = 0.6             ckappad = 0.6
+cgbo    = 0               cgbl    = 0
************************************************************
*                       temperature                        *
************************************************************
+tbgasub = 0.000473        tbgbsub = 636             kt1     = 0               kt1l    = 0
+ute     = -1.2            utl     = 0               ua1     = 0.001032        ud1     = 0
+ucste   = -0.004775       at      = 0.001           ptwgt   = 0.004           tmexp   = 0
+prt     = 0               tgidl   = -0.007          igt     = 2.5
************************************************************
*                          noise                           *
************************************************************
**)
.control
pre_osdi ~/ASAP7_FinFET_Inverter_Characterization/Xschem_ASAP7/bsimcmg_arch64.osdi
.endc



.subckt asap_7nm_nfet S G D B l=7e-009 nfin=13
	nnmos_finfet S G D B BSIMCMG_osdi_N l=7e-009 nfin=13
.ends asap_7nm_nfet

.model BSIMCMG_osdi_N BSIMCMG_va (
+ TYPE = 1
************************************************************
*                         general                          *
************************************************************
+version = 107             bulkmod = 1               igcmod  = 1               igbmod  = 0
+gidlmod = 1               iimod   = 0               geomod  = 1               rdsmod  = 0
+rgatemod= 0               rgeomod = 0               shmod   = 0               nqsmod  = 0
+coremod = 0               cgeomod = 0               capmod  = 0               tnom    = 25
+eot     = 1e-009          eotbox  = 1.4e-007        eotacc  = 1e-010          tfin    = 6.5e-009
+toxp    = 2.1e-009        nbody   = 1e+022          phig    = 4.2466          epsrox  = 3.9
+epsrsub = 11.9            easub   = 4.05            ni0sub  = 1.1e+016        bg0sub  = 1.17
+nc0sub  = 2.86e+025       nsd     = 2e+026          ngate   = 0               nseg    = 5
+l       = 2.1e-008        xl      = 1e-009          lint    = -2e-009         dlc     = 0
+dlbin   = 0               hfin    = 3.2e-008        deltaw  = 0               deltawcv= 0
+sdterm  = 0               epsrsp  = 3.9             nfin    = 1
+toxg    = 1.80e-009
************************************************************
*                            dc                            *
************************************************************
+cit     = 0               cdsc    = 0.01            cdscd   = 0.01            dvt0    = 0.05
+dvt1    = 0.47            phin    = 0.05            eta0    = 0.07            dsub    = 0.35
+k1rsce  = 0               lpe0    = 0               dvtshift= 0               qmfactor= 2.5
+etaqm   = 0.54            qm0     = 0.001           pqm     = 0.66            u0      = 0.0303
+etamob  = 2               up      = 0               ua      = 0.55            eu      = 1.2
+ud      = 0               ucs     = 1               rdswmin = 0               rdsw    = 200
+wr      = 1               rswmin  = 0               rdwmin  = 0               rshs    = 0
+rshd    = 0               vsat    = 70000           deltavsat= 0.2             ksativ  = 2
+mexp    = 4               ptwg    = 30              pclm    = 0.05            pclmg   = 0
+pdibl1  = 0               pdibl2  = 0.002           drout   = 1               pvag    = 0
+fpitch  = 2.7e-008        rth0    = 0.225           cth0    = 1.243e-006      wth0    = 2.6e-007
+lcdscd  = 5e-005          lcdscdr = 5e-005          lrdsw   = 0.2             lvsat   = 0
************************************************************
*                         leakage                          *
************************************************************
+aigc    = 0.014           bigc    = 0.005           cigc    = 0.25            dlcigs  = 1e-009
+dlcigd  = 1e-009          aigs    = 0.0115          aigd    = 0.0115          bigs    = 0.00332
+bigd    = 0.00332         cigs    = 0.35            cigd    = 0.35            poxedge = 1.1
+agidl   = 1e-012          agisl   = 1e-012          bgidl   = 10000000        bgisl   = 10000000
+egidl   = 0.35            egisl   = 0.35
************************************************************
*                            rf                            *
************************************************************
************************************************************
*                         junction                         *
************************************************************
************************************************************
*                       capacitance                        *
************************************************************
+cfs     = 0               cfd     = 0               cgso    = 1.6e-010        cgdo    = 1.6e-010
+cgsl    = 0               cgdl    = 0               ckappas = 0.6             ckappad = 0.6
+cgbo    = 0               cgbl    = 0
************************************************************
*                       temperature                        *
************************************************************
+tbgasub = 0.000473        tbgbsub = 636             kt1     = 0               kt1l    = 0
+ute     = -0.7            utl     = 0               ua1     = 0.001032        ud1     = 0
+ucste   = -0.004775       at      = 0.001           ptwgt   = 0.004           tmexp   = 0
+prt     = 0               tgidl   = -0.007          igt     = 2.5
************************************************************
*                          noise                           *
************************************************************
**)
.control
pre_osdi ~/ASAP7_FinFET_Inverter_Characterization/Xschem_ASAP7/bsimcmg_arch64.osdi
.endc


**** end user architecture code
.end
